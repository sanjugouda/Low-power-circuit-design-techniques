magic
tech scmos
timestamp 1681826354
<< polysilicon >>
rect 57 34 58 38
rect 119 34 120 38
rect 182 34 183 38
rect 245 34 246 38
rect 307 34 308 38
rect 11 30 13 32
rect 26 31 40 33
rect 26 28 28 31
rect 38 30 40 31
rect 46 30 48 32
rect 27 24 28 28
rect 11 21 13 22
rect 11 19 22 21
rect 26 20 28 24
rect 38 20 40 22
rect 46 21 48 22
rect 4 15 13 16
rect 43 19 48 21
rect 56 20 58 34
rect 73 30 75 32
rect 88 31 102 33
rect 88 28 90 31
rect 100 30 102 31
rect 108 30 110 32
rect 89 24 90 28
rect 50 18 58 20
rect 73 21 75 22
rect 73 19 84 21
rect 88 20 90 24
rect 100 20 102 22
rect 108 21 110 22
rect 0 14 13 15
rect 11 12 13 14
rect 26 12 28 14
rect 38 12 40 14
rect 50 12 52 18
rect 66 15 75 16
rect 105 19 110 21
rect 118 20 120 34
rect 136 30 138 32
rect 151 31 165 33
rect 151 28 153 31
rect 163 30 165 31
rect 171 30 173 32
rect 152 24 153 28
rect 112 18 120 20
rect 136 21 138 22
rect 136 19 147 21
rect 151 20 153 24
rect 163 20 165 22
rect 171 21 173 22
rect 62 14 75 15
rect 73 12 75 14
rect 88 12 90 14
rect 100 12 102 14
rect 112 12 114 18
rect 129 15 138 16
rect 168 19 173 21
rect 181 20 183 34
rect 199 30 201 32
rect 214 31 228 33
rect 214 28 216 31
rect 226 30 228 31
rect 234 30 236 32
rect 215 24 216 28
rect 175 18 183 20
rect 199 21 201 22
rect 199 19 210 21
rect 214 20 216 24
rect 226 20 228 22
rect 234 21 236 22
rect 125 14 138 15
rect 136 12 138 14
rect 151 12 153 14
rect 163 12 165 14
rect 175 12 177 18
rect 192 15 201 16
rect 231 19 236 21
rect 244 20 246 34
rect 261 30 263 32
rect 276 31 290 33
rect 276 28 278 31
rect 288 30 290 31
rect 296 30 298 32
rect 277 24 278 28
rect 238 18 246 20
rect 261 21 263 22
rect 261 19 272 21
rect 276 20 278 24
rect 288 20 290 22
rect 296 21 298 22
rect 188 14 201 15
rect 199 12 201 14
rect 214 12 216 14
rect 226 12 228 14
rect 238 12 240 18
rect 254 15 263 16
rect 293 19 298 21
rect 306 20 308 34
rect 300 18 308 20
rect 250 14 263 15
rect 261 12 263 14
rect 276 12 278 14
rect 288 12 290 14
rect 300 12 302 18
rect 27 8 28 12
rect 89 8 90 12
rect 152 8 153 12
rect 215 8 216 12
rect 277 8 278 12
rect 11 6 13 8
rect 26 7 28 8
rect 38 7 40 8
rect 26 5 40 7
rect 50 6 52 8
rect 73 6 75 8
rect 88 7 90 8
rect 100 7 102 8
rect 88 5 102 7
rect 112 6 114 8
rect 136 6 138 8
rect 151 7 153 8
rect 163 7 165 8
rect 151 5 165 7
rect 175 6 177 8
rect 199 6 201 8
rect 214 7 216 8
rect 226 7 228 8
rect 214 5 228 7
rect 238 6 240 8
rect 261 6 263 8
rect 276 7 278 8
rect 288 7 290 8
rect 276 5 290 7
rect 300 6 302 8
<< ndiffusion >>
rect 5 8 6 12
rect 10 8 11 12
rect 13 8 14 12
rect 18 8 19 12
rect 32 8 33 12
rect 37 8 38 12
rect 40 8 41 12
rect 45 8 50 12
rect 52 8 53 12
rect 57 8 58 12
rect 67 8 68 12
rect 72 8 73 12
rect 75 8 76 12
rect 80 8 81 12
rect 94 8 95 12
rect 99 8 100 12
rect 102 8 103 12
rect 107 8 112 12
rect 114 8 115 12
rect 119 8 120 12
rect 130 8 131 12
rect 135 8 136 12
rect 138 8 139 12
rect 143 8 144 12
rect 157 8 158 12
rect 162 8 163 12
rect 165 8 166 12
rect 170 8 175 12
rect 177 8 178 12
rect 182 8 183 12
rect 193 8 194 12
rect 198 8 199 12
rect 201 8 202 12
rect 206 8 207 12
rect 220 8 221 12
rect 225 8 226 12
rect 228 8 229 12
rect 233 8 238 12
rect 240 8 241 12
rect 245 8 246 12
rect 255 8 256 12
rect 260 8 261 12
rect 263 8 264 12
rect 268 8 269 12
rect 282 8 283 12
rect 287 8 288 12
rect 290 8 291 12
rect 295 8 300 12
rect 302 8 303 12
rect 307 8 308 12
<< pdiffusion >>
rect 5 28 11 30
rect 5 24 6 28
rect 10 24 11 28
rect 5 22 11 24
rect 13 28 19 30
rect 13 24 14 28
rect 18 24 19 28
rect 13 22 19 24
rect 32 28 38 30
rect 32 24 33 28
rect 37 24 38 28
rect 32 22 38 24
rect 40 28 46 30
rect 40 24 41 28
rect 45 24 46 28
rect 40 22 46 24
rect 48 28 54 30
rect 48 24 49 28
rect 53 24 54 28
rect 48 22 54 24
rect 67 28 73 30
rect 67 24 68 28
rect 72 24 73 28
rect 67 22 73 24
rect 75 28 81 30
rect 75 24 76 28
rect 80 24 81 28
rect 75 22 81 24
rect 94 28 100 30
rect 94 24 95 28
rect 99 24 100 28
rect 94 22 100 24
rect 102 28 108 30
rect 102 24 103 28
rect 107 24 108 28
rect 102 22 108 24
rect 110 28 116 30
rect 110 24 111 28
rect 115 24 116 28
rect 110 22 116 24
rect 130 28 136 30
rect 130 24 131 28
rect 135 24 136 28
rect 130 22 136 24
rect 138 28 144 30
rect 138 24 139 28
rect 143 24 144 28
rect 138 22 144 24
rect 157 28 163 30
rect 157 24 158 28
rect 162 24 163 28
rect 157 22 163 24
rect 165 28 171 30
rect 165 24 166 28
rect 170 24 171 28
rect 165 22 171 24
rect 173 28 179 30
rect 173 24 174 28
rect 178 24 179 28
rect 173 22 179 24
rect 193 28 199 30
rect 193 24 194 28
rect 198 24 199 28
rect 193 22 199 24
rect 201 28 207 30
rect 201 24 202 28
rect 206 24 207 28
rect 201 22 207 24
rect 220 28 226 30
rect 220 24 221 28
rect 225 24 226 28
rect 220 22 226 24
rect 228 28 234 30
rect 228 24 229 28
rect 233 24 234 28
rect 228 22 234 24
rect 236 28 242 30
rect 236 24 237 28
rect 241 24 242 28
rect 236 22 242 24
rect 255 28 261 30
rect 255 24 256 28
rect 260 24 261 28
rect 255 22 261 24
rect 263 28 269 30
rect 263 24 264 28
rect 268 24 269 28
rect 263 22 269 24
rect 282 28 288 30
rect 282 24 283 28
rect 287 24 288 28
rect 282 22 288 24
rect 290 28 296 30
rect 290 24 291 28
rect 295 24 296 28
rect 290 22 296 24
rect 298 28 304 30
rect 298 24 299 28
rect 303 24 304 28
rect 298 22 304 24
<< metal1 >>
rect 37 41 41 45
rect 45 41 95 45
rect 99 41 103 45
rect 107 41 158 45
rect 162 41 166 45
rect 170 41 221 45
rect 225 41 229 45
rect 233 41 283 45
rect 287 41 291 45
rect 295 41 309 45
rect 0 34 23 37
rect 0 19 3 34
rect 19 28 23 34
rect 33 28 37 41
rect 18 24 23 28
rect 41 34 53 38
rect 62 34 85 37
rect 41 28 45 34
rect 7 12 10 24
rect 18 12 22 15
rect 41 15 43 19
rect 50 17 53 24
rect 62 19 65 34
rect 81 28 85 34
rect 95 28 99 41
rect 80 24 85 28
rect 103 34 115 38
rect 125 34 148 37
rect 103 28 107 34
rect 41 12 45 15
rect 50 14 57 17
rect 18 8 23 12
rect 53 12 57 14
rect 69 12 72 24
rect 80 12 84 15
rect 103 15 105 19
rect 112 17 115 24
rect 125 19 128 34
rect 144 28 148 34
rect 158 28 162 41
rect 143 24 148 28
rect 166 34 178 38
rect 188 34 211 37
rect 166 28 170 34
rect 103 12 107 15
rect 112 14 119 17
rect 57 8 68 12
rect 80 8 85 12
rect 115 12 119 14
rect 132 12 135 24
rect 143 12 147 15
rect 166 15 168 19
rect 175 17 178 24
rect 188 19 191 34
rect 207 28 211 34
rect 221 28 225 41
rect 206 24 211 28
rect 229 34 241 38
rect 250 34 273 37
rect 229 28 233 34
rect 166 12 170 15
rect 175 14 182 17
rect 119 8 131 12
rect 143 8 148 12
rect 178 12 182 14
rect 195 12 198 24
rect 206 12 210 15
rect 229 15 231 19
rect 238 17 241 24
rect 250 19 253 34
rect 269 28 273 34
rect 283 28 287 41
rect 268 24 273 28
rect 291 34 303 38
rect 291 28 295 34
rect 229 12 233 15
rect 238 14 245 17
rect 206 8 211 12
rect 241 12 245 14
rect 257 12 260 24
rect 268 12 272 15
rect 291 15 293 19
rect 300 17 303 24
rect 291 12 295 15
rect 300 14 307 17
rect 245 8 256 12
rect 268 8 273 12
rect 303 12 307 14
rect 307 8 308 12
rect 33 4 37 8
rect 95 4 99 8
rect 158 4 162 8
rect 221 4 225 8
rect 283 4 287 8
rect 32 0 33 4
rect 37 0 41 4
rect 45 0 95 4
rect 99 0 103 4
rect 107 0 158 4
rect 162 0 166 4
rect 170 0 221 4
rect 225 0 229 4
rect 233 0 283 4
rect 287 0 291 4
rect 295 0 308 4
<< ntransistor >>
rect 11 8 13 12
rect 38 8 40 12
rect 50 8 52 12
rect 73 8 75 12
rect 100 8 102 12
rect 112 8 114 12
rect 136 8 138 12
rect 163 8 165 12
rect 175 8 177 12
rect 199 8 201 12
rect 226 8 228 12
rect 238 8 240 12
rect 261 8 263 12
rect 288 8 290 12
rect 300 8 302 12
<< ptransistor >>
rect 11 22 13 30
rect 38 22 40 30
rect 46 22 48 30
rect 73 22 75 30
rect 100 22 102 30
rect 108 22 110 30
rect 136 22 138 30
rect 163 22 165 30
rect 171 22 173 30
rect 199 22 201 30
rect 226 22 228 30
rect 234 22 236 30
rect 261 22 263 30
rect 288 22 290 30
rect 296 22 298 30
<< polycontact >>
rect 53 34 57 38
rect 115 34 119 38
rect 178 34 182 38
rect 241 34 245 38
rect 303 34 307 38
rect 23 24 27 28
rect 0 15 4 19
rect 18 15 22 19
rect 85 24 89 28
rect 43 15 47 19
rect 62 15 66 19
rect 80 15 84 19
rect 148 24 152 28
rect 105 15 109 19
rect 125 15 129 19
rect 143 15 147 19
rect 211 24 215 28
rect 168 15 172 19
rect 188 15 192 19
rect 206 15 210 19
rect 273 24 277 28
rect 231 15 235 19
rect 250 15 254 19
rect 268 15 272 19
rect 293 15 297 19
rect 23 8 27 12
rect 85 8 89 12
rect 148 8 152 12
rect 211 8 215 12
rect 273 8 277 12
<< ndcontact >>
rect 6 8 10 12
rect 14 8 18 12
rect 33 8 37 12
rect 41 8 45 12
rect 53 8 57 12
rect 68 8 72 12
rect 76 8 80 12
rect 95 8 99 12
rect 103 8 107 12
rect 115 8 119 12
rect 131 8 135 12
rect 139 8 143 12
rect 158 8 162 12
rect 166 8 170 12
rect 178 8 182 12
rect 194 8 198 12
rect 202 8 206 12
rect 221 8 225 12
rect 229 8 233 12
rect 241 8 245 12
rect 256 8 260 12
rect 264 8 268 12
rect 283 8 287 12
rect 291 8 295 12
rect 303 8 307 12
<< pdcontact >>
rect 6 24 10 28
rect 14 24 18 28
rect 33 24 37 28
rect 41 24 45 28
rect 49 24 53 28
rect 68 24 72 28
rect 76 24 80 28
rect 95 24 99 28
rect 103 24 107 28
rect 111 24 115 28
rect 131 24 135 28
rect 139 24 143 28
rect 158 24 162 28
rect 166 24 170 28
rect 174 24 178 28
rect 194 24 198 28
rect 202 24 206 28
rect 221 24 225 28
rect 229 24 233 28
rect 237 24 241 28
rect 256 24 260 28
rect 264 24 268 28
rect 283 24 287 28
rect 291 24 295 28
rect 299 24 303 28
<< psubstratepcontact >>
rect 33 0 37 4
rect 41 0 45 4
rect 95 0 99 4
rect 103 0 107 4
rect 158 0 162 4
rect 166 0 170 4
rect 221 0 225 4
rect 229 0 233 4
rect 283 0 287 4
rect 291 0 295 4
<< nsubstratencontact >>
rect 33 41 37 45
rect 41 41 45 45
rect 95 41 99 45
rect 103 41 107 45
rect 158 41 162 45
rect 166 41 170 45
rect 221 41 225 45
rect 229 41 233 45
rect 283 41 287 45
rect 291 41 295 45
<< labels >>
rlabel metal1 39 2 39 2 1 GND
rlabel metal1 21 26 21 26 1 GP
rlabel metal1 21 10 21 10 1 GN
rlabel metal1 9 19 9 19 1 in
rlabel metal1 40 42 40 42 5 vdd
rlabel metal1 55 15 55 15 7 out
rlabel metal1 101 2 101 2 1 GND
rlabel metal1 83 26 83 26 1 GP
rlabel metal1 83 10 83 10 1 GN
rlabel metal1 71 19 71 19 1 in
rlabel metal1 102 42 102 42 5 vdd
rlabel metal1 117 15 117 15 7 out
rlabel metal1 164 2 164 2 1 GND
rlabel metal1 146 26 146 26 1 GP
rlabel metal1 146 10 146 10 1 GN
rlabel metal1 134 19 134 19 1 in
rlabel metal1 165 42 165 42 5 vdd
rlabel metal1 180 15 180 15 7 out
rlabel metal1 227 2 227 2 1 GND
rlabel metal1 209 26 209 26 1 GP
rlabel metal1 209 10 209 10 1 GN
rlabel metal1 197 19 197 19 1 in
rlabel metal1 228 42 228 42 5 vdd
rlabel metal1 243 15 243 15 7 out
rlabel metal1 289 2 289 2 1 GND
rlabel metal1 271 26 271 26 1 GP
rlabel metal1 271 10 271 10 1 GN
rlabel metal1 259 19 259 19 1 in
rlabel metal1 290 42 290 42 5 vdd
rlabel metal1 305 15 305 15 7 out
<< end >>
